module not_gate(in, out);
	input in;
	output out;
	not(out, in);
endmodule
